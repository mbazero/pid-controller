function integer log2;
    input integer value;
    begin
        value = value-1;
        for (log2 = 0; value > 0; log2 = log2 + 1) begin
            value = value >> 1;
        end
    end
endfunction
