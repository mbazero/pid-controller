`timescale 1ns / 1ps

// pid_core -- mba 2014
// -----------------------------------------------------------
// Computes PID sum using discrete form of PID equation.
// -----------------------------------------------------------

// TODO
// - add option to set push direction

module pid_core #(
	// parameters
	parameter W_IN				= 18,								// input data width
	parameter W_OUT			= 64,								// output data width (set to be large to avoid overflow issues)
	parameter W_EP				= 16,								// width of opal kelly endpoints
	parameter COMP_LATENCY	= 1								// pid computation latency in clock cycles
	)(
	// inputs <- top level entity
	input wire									clk_in,			// system clock
	input wire									reset_in,		// system reset

	// inputs <- oversample filter
	input wire signed 	[W_IN-1:0]		data_in, 		// unsigned input data
	input wire									data_valid_in,	// input data valid signal

	// inputs <- frontpanel controller
	input wire signed		[W_EP-1:0]		setpoint_in,	// lock setpoint
	input wire signed 	[W_EP-1:0]		p_coef_in,		// proportional coefficient
	input wire signed 	[W_EP-1:0]		i_coef_in,		// integral coefficient
	input wire signed 	[W_EP-1:0]		d_coef_in,		// derivative coefficient
	input wire									lock_en_in,		// lock enable

	// outputs -> source mux
	output wire signed	[W_OUT-1:0]		data_out,		// pid filter output
	output wire									data_valid_out	// output data valid signal
   );

//////////////////////////////////////////
// local parameters
//////////////////////////////////////////

localparam MAX_OUTPUT = {1'b0, {W_OUT-1{1'b1}}};
localparam MIN_OUTPUT = ~MAX_OUTPUT;

/* state parameters */
localparam 	ST_IDLE 			= 3'd0,							// module idle, wait for valid data
				ST_COMPUTE		= 3'd1,							// compute filter output
				ST_SEND			= 3'd2, 							// send filter data downstream
				ST_WRITEBACK	= 3'd3; 							// cycle complete, writeback pid sum and error

//////////////////////////////////////////
// internal structures
//////////////////////////////////////////

/* input data */
reg signed	[W_IN-1:0]		data = 0;						// active input data

/* overflow handling */
wire 								overflow;
wire signed [W_OUT-1:0]		u_cur_rail;

/* error signals */
wire signed	[W_IN:0]			e_cur;							// current error signal
reg signed	[W_IN:0]			e_prev_0 = 0;					// most recent previous error signal
reg signed	[W_IN:0]			e_prev_1 = 0;					// second most recent previous error signal

/* z-transform coefficients */
wire signed	[W_EP+1:0]		k1, k2, k3; 					// z-transform coefficients for discrete PID filter

/* control variable (u) cur, prev, and delta vals */
reg signed	[W_OUT-1:0]		u_prev = 0;						// previous pid filter output
wire signed	[W_OUT-1:0]		u_cur; 							// current pid filter output
wire signed	[W_OUT-1:0]		delta_u;							// difference between current and previous pid filter outputs

/* state registers */
reg			[7:0] 			counter = 0; 					// intrastate counter
reg			[2:0] 			cur_state = ST_IDLE;			// current state
reg			[2:0] 			next_state = ST_IDLE; 		// next state

//////////////////////////////////////////
// combinational logic
//////////////////////////////////////////

/* compute error */
assign e_cur				= setpoint_in - data;

/* compute z-transform coefficients */
assign k1					= p_coef_in + i_coef_in + d_coef_in;
assign k2					= -p_coef_in - (d_coef_in << 1);
assign k3					= d_coef_in;

/* compute delta u */
assign delta_u				= k1*e_cur + k2*e_prev_0 + k3*e_prev_1;

/* compute u */
assign u_cur				= delta_u + u_prev;

/* check for overflow */
assign overflow 			= (delta_u[W_OUT-1] == u_prev[W_OUT-1])
									&& (u_prev[W_OUT-1] != u_cur[W_OUT-1]);
assign u_cur_rail			= (u_prev[W_OUT-1] == 0) ? MAX_OUTPUT : MIN_OUTPUT;

/* data out */
assign data_out			= ( overflow ) ? u_cur_rail : u_cur;
assign data_valid_out	= ( cur_state == ST_SEND );

//////////////////////////////////////////
// sequential logic
//////////////////////////////////////////

/* data register */
always @ ( posedge clk_in ) begin
	if (( reset_in == 1 ) | ( lock_en_in == 0 )) begin
		data <= 0;
	end else if (( data_valid_in == 1 ) & ( cur_state == ST_IDLE )) begin
		data <= data_in;
	end
end

/* previous error and output registers */
always @( posedge clk_in ) begin
	if (( reset_in == 1 ) | ( lock_en_in == 0 )) begin
		u_prev	<= 0;
		e_prev_0	<= 0;
		e_prev_1	<= 0;
	end else if ( cur_state == ST_WRITEBACK ) begin
		u_prev	<= data_out;
		e_prev_0	<= e_cur;
		e_prev_1	<= e_prev_0;
	end
end

//////////////////////////////////////////
// state machine
//////////////////////////////////////////

/* state sequential logic */
always @( posedge clk_in ) begin
	if ( reset_in == 1 ) begin
		cur_state <= ST_IDLE;
	end else begin
		cur_state <= next_state;
	end
end

/* state counter sequential logic */
always @( posedge clk_in ) begin
	if ( reset_in == 1 ) begin
		counter <= 0;
	end else if ( cur_state != next_state ) begin
		counter <= 0;
	end else begin
		counter <= counter + 1;
	end
end

/* next state combinational logic */
always @( * ) begin
	next_state <= cur_state; // default assignment if no case and condition is satisfied
	case ( cur_state )
		ST_IDLE: begin
			if ( data_valid_in == 1 )			next_state <= ST_COMPUTE;
		end
		ST_COMPUTE: begin
			if ( counter == COMP_LATENCY-1 )	next_state <= ST_SEND;
		end
		ST_SEND: 									next_state <= ST_WRITEBACK;
		ST_WRITEBACK:								next_state <= ST_IDLE;
	endcase
end

endmodule
