parameter mask							= 32'hffffffff;
